`ifndef DATAPATH_SV
`define DATAPATH_SV

`define BAD_MUX_SEL $fatal("%0t %s %0d: Illegal mux select", $time, `__FILE__, `__LINE__)
import rv32i_types::*;

module datapath(
    input clk,
    input rst,
    // from i-cache
    input rv32i_word icache_rdata,
    // to i-cache
    output [31:0] icache_addr,
    output icache_read,
    // from d-cache
    input rv32i_word dcache_rdata,
    // to d-cache
    output [31:0] dcache_addr,
    output dcache_read,
    output dcache_write,
    output logic [3:0] dcache_byte_en,
    output rv32i_word dcache_wdata,
    // NOTE byte_en is generated by datapath
    // from control
    input rv32i_control_word ctl_word,
    // to control
    output rv32i_funct_word fd_word,
    output rv32i_funct_word de_word,
    output rv32i_funct_word em_word,
    output rv32i_funct_word mw_word
);

// internal signals
// signals between latches
logic fd_valid_out;
logic [31:0] fd_instr_latch_out, fd_pc_latch_out, fd_rs1_latch_out, fd_rs2_latch_out;
logic [31:0] fd_alu_latch_out, fd_dc_latch_out;
// logic [31:0] marmux_out;
logic [2:0] fd_funct3;
logic [6:0] fd_funct7;
rv32i_opcode fd_opcode;
logic [31:0] fd_i_imm, fd_s_imm, fd_b_imm, fd_u_imm, fd_j_imm;
logic [4:0] fd_rs1, fd_rs2, fd_rd;

logic de_valid_out;
logic [31:0] de_instr_latch_out, de_pc_latch_out, de_rs1_latch_out, de_rs2_latch_out;
logic [31:0] de_alu_latch_out, de_dc_latch_out;
logic [2:0] de_funct3;
logic [6:0] de_funct7;
rv32i_opcode de_opcode;
logic [31:0] de_i_imm, de_s_imm, de_b_imm, de_u_imm, de_j_imm;
logic [4:0] de_rs1, de_rs2, de_rd;

logic em_valid_out;
logic [31:0] em_instr_latch_out, em_pc_latch_out, em_rs1_latch_out, em_rs2_latch_out;
logic [31:0] em_alu_latch_out, em_dc_latch_out;
logic [2:0] em_funct3;
logic [6:0] em_funct7;
rv32i_opcode em_opcode;
logic [31:0] em_i_imm, em_s_imm, em_b_imm, em_u_imm, em_j_imm;
logic [4:0] em_rs1, em_rs2, em_rd;

logic mw_valid_out;
logic [31:0] mw_instr_latch_out, mw_pc_latch_out, mw_rs1_latch_out, mw_rs2_latch_out;
logic [31:0] mw_alu_latch_out, mw_dc_latch_out;
logic [2:0] mw_funct3;
logic [6:0] mw_funct7;
rv32i_opcode mw_opcode;
logic [31:0] mw_i_imm, mw_s_imm, mw_b_imm, mw_u_imm, mw_j_imm;
logic [4:0] mw_rs1, mw_rs2, mw_rd;


// IF Signals
rv32i_word pcmux_out, pc_out;
// ID signals
logic [31:0] rs1_out, rs2_out;
logic add_bubble;
// EX signals
logic br_en;
logic [31:0] cmpmux_out;
logic [31:0] alu_out;
logic [31:0] arithmux_out, alumux1_out, alumux2_out;
logic keep_delay_slot;
// MEM signals
// WB signals
logic [31:0] regfilemux_out;

// forwarder signals
logic [31:0] rs1_forwarder_out;
logic [31:0] rs2_forwarder_out;

// instantiate alu cmp regfile pc_reg
alu ALU(
    .aluop(ctl_word.aluop),
    .a(alumux1_out), .b(alumux2_out),
    .f(alu_out)
);

cmp CMP(
    .cmpop(ctl_word.cmpop),
    .a(rs1_forwarder_out), .b(cmpmux_out),
    .br_en(br_en)
);

regfile REGFILE(
    .clk(clk), .rst(rst),
    .load(ctl_word.load_regfile), .in(regfilemux_out), .dest(mw_rd),
    .src_a(fd_rs1), .reg_a(rs1_out),
    .src_b(fd_rs2), .reg_b(rs2_out)
);

pc_register PC_REGISTER(
    .clk(clk), .rst(rst),
    .load(ctl_word.load_pc & ~add_bubble), .in(pcmux_out), .out(pc_out)
);

forwarder FORWARDER(.*);


// instatiate latches between stages
// FIXME : timing of load pc and write pc to fd latch
ilatch FD_LATCH( // IF/ID latch
    .clk(clk), .rst(rst), .load(ctl_word.load_latch & ~add_bubble),
    .valid_in(1'b1), .valid_ctl(keep_delay_slot), .valid_out(fd_valid_out),
    .instr_latch_in(icache_rdata), .instr_latch_out(fd_instr_latch_out),
    .pc_latch_in(pc_out), .pc_latch_out(fd_pc_latch_out),
    .rs1_latch_in(32'b0), .rs1_latch_out(fd_rs1_latch_out),
    .rs2_latch_in(32'b0), .rs2_latch_out(fd_rs2_latch_out),
    .alu_latch_in(32'b0), .alu_latch_out(fd_alu_latch_out),
    .dc_latch_in(32'b0), .dc_latch_out(fd_dc_latch_out),
    // not passed
    .funct3(fd_funct3), .funct7(fd_funct7), .opcode(fd_opcode),
    .i_imm(fd_i_imm), .s_imm(fd_s_imm), .b_imm(fd_b_imm), .u_imm(fd_u_imm), .j_imm(fd_j_imm),
    .rs1(fd_rs1), .rs2(fd_rs2), .rd(fd_rd)
);

ilatch DE_LATCH( // ID/EX latch
    .clk(clk), .rst(rst), .load(ctl_word.load_latch),
    .valid_in(fd_valid_out), .valid_ctl(keep_delay_slot & ~add_bubble), .valid_out(de_valid_out),
    .instr_latch_in(fd_instr_latch_out), .instr_latch_out(de_instr_latch_out),
    .pc_latch_in(fd_pc_latch_out), .pc_latch_out(de_pc_latch_out),
    .rs1_latch_in(rs1_out), .rs1_latch_out(de_rs1_latch_out),
    .rs2_latch_in(rs2_out), .rs2_latch_out(de_rs2_latch_out),
    .alu_latch_in(32'b0), .alu_latch_out(de_alu_latch_out),
    .dc_latch_in(32'b0), .dc_latch_out(de_dc_latch_out),
    // not passed
    .funct3(de_funct3), .funct7(de_funct7), .opcode(de_opcode),
    .i_imm(de_i_imm), .s_imm(de_s_imm), .b_imm(de_b_imm), .u_imm(de_u_imm), .j_imm(de_j_imm),
    .rs1(de_rs1), .rs2(de_rs2), .rd(de_rd)
);

ilatch EM_LATCH( // EX/MEM latch
    .clk(clk), .rst(rst), .load(ctl_word.load_latch),
    .valid_in(de_valid_out), .valid_ctl(1'b1), .valid_out(em_valid_out),
    .instr_latch_in(de_instr_latch_out), .instr_latch_out(em_instr_latch_out),
    .pc_latch_in(de_pc_latch_out), .pc_latch_out(em_pc_latch_out),
    .rs1_latch_in(rs1_forwarder_out), .rs1_latch_out(em_rs1_latch_out),
    .rs2_latch_in(rs2_forwarder_out), .rs2_latch_out(em_rs2_latch_out),
    .alu_latch_in(arithmux_out), .alu_latch_out(em_alu_latch_out),
    .dc_latch_in(32'b0), .dc_latch_out(em_dc_latch_out),
    // not passed
    .funct3(em_funct3), .funct7(em_funct7), .opcode(em_opcode),
    .i_imm(em_i_imm), .s_imm(em_s_imm), .b_imm(em_b_imm), .u_imm(em_u_imm), .j_imm(em_j_imm),
    .rs1(em_rs1), .rs2(em_rs2), .rd(em_rd)
);

ilatch MW_LATCH( // MEM/WB latch
    .clk(clk), .rst(rst), .load(ctl_word.load_latch),
    .valid_in(em_valid_out), .valid_ctl(1'b1), .valid_out(mw_valid_out),
    .instr_latch_in(em_instr_latch_out), .instr_latch_out(mw_instr_latch_out),
    .pc_latch_in(em_pc_latch_out), .pc_latch_out(mw_pc_latch_out),
    .rs1_latch_in(em_rs1_latch_out), .rs1_latch_out(mw_rs1_latch_out),
    .rs2_latch_in(em_rs2_latch_out), .rs2_latch_out(mw_rs2_latch_out),
    .alu_latch_in(em_alu_latch_out), .alu_latch_out(mw_alu_latch_out),
    .dc_latch_in(dcache_rdata), .dc_latch_out(mw_dc_latch_out),
    // not passed
    .funct3(mw_funct3), .funct7(mw_funct7), .opcode(mw_opcode),
    .i_imm(mw_i_imm), .s_imm(mw_s_imm), .b_imm(mw_b_imm), .u_imm(mw_u_imm), .j_imm(mw_j_imm),
    .rs1(mw_rs1), .rs2(mw_rs2), .rd(mw_rd)
);

assign fd_word.funct3      = fd_funct3;
assign fd_word.funct7      = fd_funct7;
assign fd_word.opcode      = fd_opcode;
assign fd_word.word_valid  = fd_valid_out;

assign de_word.funct3      = de_funct3;
assign de_word.funct7      = de_funct7;
assign de_word.opcode      = de_opcode;
assign de_word.word_valid  = de_valid_out;

assign em_word.funct3      = em_funct3;
assign em_word.funct7      = em_funct7;
assign em_word.opcode      = em_opcode;
assign em_word.word_valid  = em_valid_out;

assign mw_word.funct3      = mw_funct3;
assign mw_word.funct7      = mw_funct7;
assign mw_word.opcode      = mw_opcode;
assign mw_word.word_valid  = mw_valid_out;
// output signal assignment
assign icache_addr = pc_out;
assign icache_read = ctl_word.icache_read;
assign dcache_addr = em_alu_latch_out;
assign dcache_read = ctl_word.dcache_read;
assign dcache_write = ctl_word.dcache_write;


function void set_default();
    pcmux_out = pc_out + 4;
    // marmux_out = pc_out;
    alumux1_out = rs1_forwarder_out;
    alumux2_out = de_i_imm;
    cmpmux_out = rs2_forwarder_out;
    arithmux_out = alu_out;
    dcache_byte_en = 4'b1111;
    dcache_wdata = em_rs2_latch_out;
    regfilemux_out = mw_alu_latch_out;
endfunction

// muxes
always_comb
begin
    // set default to prevent "not purely combinational logic"
    set_default();
    // TODO muxes for IF stage
    // iaddrmux
    // FIXME need to change marmux and pcmux to make this work
    unique case(ctl_word.iaddrmux_sel)
        iaddrmux::always_pc : begin
            pcmux_out = pc_out + 4;
            // marmux_out = pc_out;
        end
        iaddrmux::always_alu: begin
            pcmux_out = {alu_out[31:1],1'b0};
            // marmux_out = {alu_out[31:1],1'b0};
        end
        iaddrmux::br_en     : begin
            // pc_in_mux
            // NOTE: pcmux_sel/ marmux_sel = iaddrmux_out
            // NOTE last bit of alu is always ignored
            unique case (br_en)
                pcmux::pc_plus4: pcmux_out = pc_out + 4;
                pcmux::alu_plus4: pcmux_out = {alu_out[31:1],1'b0};
                default: `BAD_MUX_SEL;
            endcase
            // // mar_mux
            // unique case (br_en)
            //     marmux::pc_out: marmux_out = pc_out;
            //     marmux::alu_out: marmux_out = {alu_out[31:1],1'b0};
            //     default: `BAD_MUX_SEL;
            // endcase            
        end
        default: `BAD_MUX_SEL;
    endcase

    // TODO muxes for ID stage
    if(de_valid_out && de_opcode == op_load && de_rd != '0 &&
       (de_rd == fd_rs1 || de_rd == fd_rs2)) // FIXME what about invalid fd or de?
        add_bubble = 1'b1;
    else
        add_bubble = 1'b0; // default is not add

    // TODO muxes for EX stage
    // alu_src1_mux
    unique case(ctl_word.alumux1_sel)
        alumux::rs1_out : alumux1_out = rs1_forwarder_out;
        alumux::pc_out  : alumux1_out = de_pc_latch_out;
        default: `BAD_MUX_SEL;
    endcase
    // alu_src2_mux
    unique case(ctl_word.alumux2_sel)
        alumux::i_imm   : alumux2_out = de_i_imm;
        alumux::u_imm   : alumux2_out = de_u_imm;
        alumux::b_imm   : alumux2_out = de_b_imm;
        alumux::s_imm   : alumux2_out = de_s_imm;
        alumux::j_imm   : alumux2_out = de_j_imm;
        alumux::rs2_out : alumux2_out = rs2_forwarder_out;
        default: `BAD_MUX_SEL;
    endcase
    // cmp_src2_mux
    unique case(ctl_word.cmpmux_sel)
        cmpmux::rs2_out: cmpmux_out = rs2_forwarder_out;
        cmpmux::i_imm  : cmpmux_out = de_i_imm;
        default: `BAD_MUX_SEL;
    endcase
    // arithmux
    unique case(ctl_word.arithmux_sel)
        alumux::alu_out: arithmux_out = alu_out;
        alumux::cmp_out: arithmux_out = {31'd0, br_en};
        default: `BAD_MUX_SEL;
    endcase
    // whether to keep delay slot
    if ((ctl_word.iaddrmux_sel == iaddrmux::always_alu) || (ctl_word.iaddrmux_sel == iaddrmux::br_en && br_en))
        keep_delay_slot = 1'b0;
    else
        keep_delay_slot = 1'b1;

    // TODO muxes for MEM stage
    case(store_funct3_t'(em_funct3))
        sb: begin
            dcache_byte_en = 4'b0001 << em_alu_latch_out[1:0];
            dcache_wdata = em_rs2_latch_out << {em_alu_latch_out[1:0], 3'd0};
        end
        sh: begin
            dcache_byte_en = 4'b0011 << {em_alu_latch_out[1], 1'b0};
            dcache_wdata = em_rs2_latch_out << {em_alu_latch_out[1], 4'd0};
        end
        sw: begin
            dcache_byte_en = 4'b1111;
            dcache_wdata = em_rs2_latch_out;
        end
        default: begin
            dcache_byte_en = '0;
            dcache_wdata = '0;
        end
    endcase

    // TODO muxes for WB stage
    // regfile_in_mux
    unique case (ctl_word.regfilemux_sel)
        regfilemux::alu_out:  regfilemux_out = mw_alu_latch_out;
        // regfilemux::br_en:    regfilemux_out = br_en;
        regfilemux::u_imm:    regfilemux_out = mw_u_imm;
        regfilemux::lw:       regfilemux_out = mw_dc_latch_out;
        regfilemux::pc_plus4: regfilemux_out = mw_pc_latch_out + 4;
        regfilemux::lb:
            case(mw_alu_latch_out[1:0])
                2'b00: regfilemux_out = {{24{mw_dc_latch_out[ 7]}}, mw_dc_latch_out[ 7: 0]};
                2'b01: regfilemux_out = {{24{mw_dc_latch_out[15]}}, mw_dc_latch_out[15: 8]};
                2'b10: regfilemux_out = {{24{mw_dc_latch_out[23]}}, mw_dc_latch_out[23:16]};
                2'b11: regfilemux_out = {{24{mw_dc_latch_out[31]}}, mw_dc_latch_out[31:24]};
            endcase
        regfilemux::lbu:
            case(mw_alu_latch_out[1:0])
                2'b00: regfilemux_out = {24'd0, mw_dc_latch_out[ 7: 0]};
                2'b01: regfilemux_out = {24'd0, mw_dc_latch_out[15: 8]};
                2'b10: regfilemux_out = {24'd0, mw_dc_latch_out[23:16]};
                2'b11: regfilemux_out = {24'd0, mw_dc_latch_out[31:24]};
            endcase
        regfilemux::lh:
            case(mw_alu_latch_out[1])
                1'b0: regfilemux_out = {{16{mw_dc_latch_out[15]}}, mw_dc_latch_out[15: 0]};
                1'b1: regfilemux_out = {{16{mw_dc_latch_out[31]}}, mw_dc_latch_out[31:16]};
            endcase
        regfilemux::lhu:
            case(mw_alu_latch_out[1])
                1'b0: regfilemux_out = {16'd0, mw_dc_latch_out[15: 0]};
                1'b1: regfilemux_out = {16'd0, mw_dc_latch_out[31:16]};
            endcase
        default: `BAD_MUX_SEL;
    endcase

end

endmodule : datapath

`endif
